--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   17:54:33 05/04/2024
-- Design Name:   
-- Module Name:   /home/rahul/Desktop/13031122015/ALU_4bit/alu_test.vhd
-- Project Name:  ALU_4bit
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: alu_rtl
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY alu_test IS
END alu_test;
 
ARCHITECTURE behavior OF alu_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT alu_rtl
    PORT(
         A : IN  std_logic_vector(3 downto 0);
         B : IN  std_logic_vector(3 downto 0);
         S : IN  std_logic_vector(2 downto 0);
         ALU_Out : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal A : std_logic_vector(3 downto 0) := (others => '0');
   signal B : std_logic_vector(3 downto 0) := (others => '0');
   signal S : std_logic_vector(2 downto 0) := (others => '0');

 	--Outputs
   signal ALU_Out : std_logic_vector(3 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: alu_rtl PORT MAP (
          A => A,
          B => B,
          S => S,
          ALU_Out => ALU_Out
        );

   -- Clock process definitions
 

   -- Stimulus process
   stim_proc: process
   begin	
	A <= "0001";
	B <= "0010";
	
	S <= "000";
	wait for 1 ps;
	S <= "001";
	wait for 1 ps;
	S <= "010";
	wait for 1 ps;
	S <= "011";
	wait for 1 ps;
	S <= "100";
	wait for 1 ps;
	S <= "101";
	wait for 1 ps;
	S <= "110";
	wait for 1 ps;
	S <= "111";
	wait for 1 ps;
	
	
   end process;

END;
